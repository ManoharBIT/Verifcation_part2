// apb_pkg.sv

package apb_pkg; 
  // apb agent files
  `include "apb_xtn.sv"
  `include "apb_sequencer.sv"
  `include "apb_agent_config.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_agent.sv"
  `include "apb_env_config.sv"
  `include "apb_sb.sv"
  `include "apb_env.sv"
endpackage