//interface

interface intf();
  
  logic a;
  logic b;
  logic c;
  logic sum;
  logic carry;
  
  //clocking block
  //modport
  
endinterface/*interface fa_if(input logic clk);
    logic a, b, cin;
    logic sum, cout;
endinterface
*/ 